// This is a model of TSV

module TSV(input i, output o);
  assign o = i;
endmodule
